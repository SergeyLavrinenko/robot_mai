/* Definition of the `ping` component. */

component echo.Configuration

endpoints {
    /* Declaration of a named implementation of the "Ping" interface. */
    getConfiguration : echo.Configuration
}
